PK   :�W8x �  �<    cirkitFile.json�]m��6��+���(����..��2@�3C����=v�۝I.��~�$�-��ʪrOv$�X,����C�[�[m��j�[ux��w�{���Oš�R\~ʖ���nuܯ~=�����'�?�d�����U��ʰR!ER�U�(�.�<MYb2��M�x��+���q9�9�5���\�k\�����g��96X�!qǑ��y�֙2����D�R%�ެ���dR��Ȅ�E�����U���u��LXU�D�9O
%�$���ް��<��ӵ�t]�ņ�<O��m��z���I���Ne��Fv�\-�\8r�p�,2�eQ���y��I����'l�n
a6EU��zL�շ���8W%3E��Yf[�,)6��G�B�Z��zd{5���y�%@����y|{5�oO���j_o����j_m0�`a�����k�DGB�#�װ�K���*��޺�����2+�D��V�7�Z�,���&/��2[1� �=��f�2_��G�_ �/���D�@�_ �/��H�H�
$�
$�$�?������H��8�@Ǔ�����[q7�l�U��:D��V�:^1T�<>���f�c_t����r�γ���]�v�.�$ϔJ*i*;w�L��6F��Ҡ�c�aP�1��z��@=���c��s,��Yaz��=@=���bz�-hP��s���9��t�z�1=�(&A�Ǳ��P<�QD�QL����FqY4���f�(.�o���q��D��!pX�4���;��o	s7p��Ot���ظ�4L��s���!��-�CD�1R����c�t=�<<�{��9F�@��s�H��!�瘇t1L���ñ��P<���!�o�E=<�����fQ���%��S �7`�P�A���a��� V�n�g�6���ۀ������m�j`���6`50/�z���Jp�X��G����%5\oV�2#������3H��)	�ϕ^��+�l�%�̰ϗ^��+��9�fؠ��T�s}�zܸy1�Y�#������an�1�:r�	R�0���6�ݻ�����|b�k��m��A�E�h�$Z�M�%%�bH�d$Zr�������ů���¨i \mʚ�u��/EaN�aNbN�bѠ8�d)�5�������O.)�;Z&�-����-��	����ɥ}w�uD�A��~ ~��B�9���@�0jh0���ذf��łł��iP,hP,hP,hP,h�XРX�P��A��A��A�$r%hP,iP,'Q}��@�"t��g�K	�t}�`�A_??A���eu���J����6y�	۵����4��z�L��o�-$S�#�gh��⻜�l9�A�֝-\+��b�S\.Q��l�fL-�N�k�����W�45-�TjSDb���k;4�]L�>EiK#Ή^|��T(k�(M�D^b�L�3����H8�x<.N#������4�w�ȡ)��DM�'rh��8�C�`ǉ��:N����q"����94mt�ȡ)��DN�'rpf�8���,ǉ�/9N����q"g1�94!q�������Y9��meV� �"�O�J��(r@��FHcQ�;+��ƢȱyV�!�E����C�".ܬ�C�"ѭYɈ4Ee�Ri,���f%*1$iSibы�yI�D6�7�&�2���HdySi:y[��p^ �&����v���1�t,�6clW=�&y�D� �"I�(-�DKJ�Őh�H��4�#/z9|9~9�9�9�9�9�9���$��cx-4�L.(p�^��rg��L.&p�^��Rg����4���cjh <��3���`xz?�g�����A�bA�bA�bA�bA�bA�bA�bA�bI�bI�bI�JРXҠXN��1��29O��1���Yg��L�8c��Ɩ�9g��L.$p�^��f ��k��
�c�#/z��rx�� O{���154����c�7�bp�^��R g��L.p�^��2 g��L.p�^���g���A�4��3��� x���cx-�y��1F��S)�輌1�"h��1FbQda��#�(���e��XY��2�H,�l^�2�H,�l��2�H,�l��2�H,�l��2�h����4�=��c46�7���O33c��&2����ff���DF�=M_��?��V���Ž��ŗ�zZ=>��\mw����������(g��Uku�@��z������P�9LߘwIsTϘ2��g̛��3�@c���F6fea^�S��y�5�d���~�%��%Lϸ�
(��@�G1ݣ�E��#
�9(D���a�ܙ?�@Xcyf��oZ+�=C��v�6�=�N�F�zv�o.�}�/Lt�Q��b�A�F��sn|�f� ��:S�D�7cYhu���S������Ӌ]:���vZ������a���A�Q^'�7����L�@(� �x��
�RDF-�#�^�@�0�����h����	���+��0�	�hH��o�1� 6r��$h���&��7���XA2#�p��c��t,����4�sS#����}�U<��J�gԂW	��t� G}\�����ݝ�������B�������YaF�^ �Kd{�l���Sd{�l�!��X���E �B�I�c�?IĞ>�����h�Y�-Ǣ�caۼ���ë��a~�hdU��`ڏ�)p�L�Z���Y"��<��#\��4 ��ux��,9�SX%���A��E�k�%wP<�ũ@3%��S�ũ��T`�R`�)��)�H�X$J,%z��"Qb�(G�.��ip�"���;Y����\!�e��r`�p͜�u�0���n8=u�����bn�(�dU�P�ɑ�ԏA_&��8s[���0�H��e�YxY��>�����.�����94i�n��{�P�K#��z�� ԏ�\~������mb��>}rW��C�&��p͟�:L� |�W꫋m;�r@u���o;�Au�u�4P�I��o;��A}�e�v�Մ�Pɴ�m^_h`j>�����@]d��K&��W�V���a�y��Vx��yU��Vx��y���Vx�yՄ�Vxa�y��Vx�㼪AH+�P޼JAH+�x��@H+��⼊@X�" O���Y�k��u����
?X;H�#���H��U��K���~<�_���k[�d1�Ǔ���$,��/����`�Z;wݹ��Mtw�qv��hN}�I�9�6'��?m�����/�`��5��/ ���1��˵��p-�k!\�Z�B�ҵ���l�q-�k!��H4��J.�(ih@b7<k��Ae��r��'������n��C��;����W�c���Ƙ������R�,?:�0[Eˏ� ����Zc������l�-?�0[�ˏ�"�7�H�EF��n�!G�-��G�1��a��1(���㡘�	]��b�A����0�+��W�s������=�_���'&c	uw��2�d�S�c�������cQW☜0o(El�}�"S~�[ؚש;姤��y�w_αGW���XW�8������qKl��w���Ht���Hv���Hu���Hw���(���#�=2���{�����Q�=����p��p���O��������ӈpH�iH�?&�4&�~�
?�
��������"N�"�q�q���3N�1�������a�tt�D�z��r�T�'��*)�:�k��ʴ9�r�ʕX���Z%���2��d�]��t�P�Gk���U���ᩲ,i����ݪ����z^�O+����g�ѻ���:�U|���s�q`G��x��~��gW|vwO��ߊ�g�7Kdn�w[k����ӧ���v�f�.�kg�}�T~�>m����C�?��CU.�vd�4}.v�u�9>\��x�b/f��,������v�kc�	�*k���i{��퀼�)�c"7*U��%7�[6��;��r��Jd�%M!�f�tbg�n�E)EU(f�*k�v�t,v��(�\����ְE���d�=l�n^�+s����}�������k����k���i��l�����2�wc���8s�8K;u&��	�ș�3�V��4�>�&�9�Ns;a�~׭\�k����ڏ��}ݼ5/��g��UgN��ԥ�:q�a9ݎrv2/"&�p2�r����|�|L�|��<����x�YW��>>���/��]t���1��`	��s���m�r�T�<��|�4�ݩ���%m��ԕX�I��*�,��rb���Ȕʳ!m�n膴iw�!i��n�;�df�
�t��Խ�_D�4��0mY_����"f8�6#@���&#bZ��̶�-c m}�L��:�:ۡ:�> ' �M@* ��T 5� h|�fR���	H �
�% ��/BK@* ��T +�0�|���%�"b�ݥ��u[�eyPY@*�K
����������U���-���b����$��A����g�4�Lj!eR�sE��1�=�dM�Ho%� vP�V�R��������O�~"O2�6��<��/	�R�7 ����?��#Ǎqǁ��~����V��)���&��2IE�����^mri�=�h#�� FZ��vLg�%\��T��Ͻ����� �Dn�[�cm�-���[j��á��u��:/ڞ0�u����R���t#�!@�]�X�%���bO����D��T��B�D�\b��M�������7M쑽ۋ�MD�6a]q~�5MXn��WwT���-��ka�OZ�S�����]tm��6-��ӗ|1��m����OLۆg�y�6a��ڗ�i!O,l��Xʻ4\�����T	�:���ug���N_���`��e&=�MD�:ji�qލ�A�R�sfq5PܞS���3bѕڙq�i�X��-�	��~�<��uV�'U��[Gm��δNʂ��Ϊ�}ѮG-�dM�N��R�3���E]>�����8=y���b-ҋޅ����D��!bO�����'<���na��ep��h�L���~��������9j�Y��+��þ(�ס�ɬ/�S�u�ƺ"���kSIn��u����u���*1���r0c���jq����-k��ڿNͼ���?��fƏ�G��;p�N�۰�E�Dny�)�|ٖ�ON����S������]ֵ�}��K���b�*�?ߖ�;T���l�/��~��]���a���������w��H����Cq8���~(�G�s�mծ�L�nt�/?�g��о��vw|W?5�������]P�T�s~nٓ�����wK=g�YY>��8�eHL����؋�v����W��>@򊱬"� �������^�,��Xt�{�1\V�M�I�	©�i�g���D2��|�X���[2� a� a� a� a� "@2��|�D2ӵ�)���#'�GN��|8$�=$�=z�����Ҳ�GF��)8�y��0��0�����bЭ%��G	CCC
3)�9Rs���p1�µR��H����#%G:�92s���b�m��l�����&�&����9�9z7Tp1(s�r�)��������H��f����@,6���M�i��tC	)u��6\:/Zڿ���C����2GQ�:���R�X)m�t^�����C�#.��E����6yM�"pQǷh�[�f]�(AЬ��j�X�Y��n�aM�&mPs^L���u�#��b}��BL0�oF���bQ��	�0pu]���J�п��.��p�<��a��KaWz�ܵ�+��4��D^���t̩�ǜ�|���_�#�P7�0j�C���ix�d)��`�B�\���82��
̟�!m���r���ЁP��ŀ���&��_������Z��zɵ`�S�,_umT!I� �����5Ƒ-�Y�W,�Bat'�)����{�ŀ@�{��ghs
`�`mN=�)���L��׉�n�T�r�ng�����"�o��g\�yʗz+~u���6x����+'�k�s91�A)��~*�/����WwS��#�W�z-R2RRy��������uӰ�����ME��Y�OA��B�2$�T�P9n
Iq��!.�Xĉ��{�.ص�9o�&���W�z��AKb ł�2l��fߌ?9*�Z���
��>���Z��@6d�؁��Nva�5�f�/U�)xK{d���"8C��Ȧi�lip��l��[���t���l���#[x��	��7����7�^�c֬,��*<�C���� ��1K�:f}K@���Q���Y��PH��t�C��K�b��v��.Bz�C�b��Qa�Q��"�M +oO|O&�¼Y;�+X����A�R�+��0�@�!�T�RΑ�� �����a/���#P�����ԩ�T
zx�YCs���@�c\�>z�mTnŬ�їѣKi v'�T�6@�R1��`X*r�]e9��u��ij0�s��0�Z0vƳ@0�"�=��¤�]9L�Iy�����.
"� �J�l~�,��a[<<-�����l��*,v������?��On�?~]|�?PK
   :�W8x �  �<                  cirkitFile.jsonPK      =   =    